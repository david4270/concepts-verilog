

module proc();

endmodule