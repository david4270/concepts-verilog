`timescale 1ns/1ns
`include "proc.sv"

module proc_tb();
    
endmodule